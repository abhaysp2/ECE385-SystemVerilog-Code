// lab7_soc_subsystemA_0.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module lab7_soc_subsystemA_0 (
	);

endmodule
